library IEEE;
use IEEE.std_logic_1164.all;

entity comparator_33000 is 
    port (
        

    );
    end;

architecture comparator_33000_arch of comparator_33000 is
end;