library IEEE;
use IEEE.std_logic_1164.all;

entity comparator_33000 is 
    port (
        A : in std_logic_vector(21 downto 0);
        B : in std_logic_vector(21 downto 0);
        q : out std_logic
    );
    end;

architecture comparator_33000_arch of comparator_33000 is
end;