library IEEE;
use IEEE.std_logic_1164.all;

entity binary_counter is
    port (
        clk : in std_logic;
        q_reg : out std_logic;
        q_BCD : out std_logic; 
    );
    end;

architecture binary_counter_arch of binary_counter is
end;